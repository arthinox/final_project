module keyboard_ctrl {
	input [7:0] keycode,
	output 
};

// Code that takes keyboard input and converts into data used by waveform generator

always_comb
	begin
		case (keycode)
		
	end

endmodule
