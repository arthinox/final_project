module i2s (
	input I2S_MCLK, I2S_DIN,
	output I2S_LRCLK, I2S_SCLK,
	output I2S_DOUT
);


endmodule
