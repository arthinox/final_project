module wave_generator (
	input CLK, Reset,
	input [2:0] tone,
	output [23:0] sample
);

	
endmodule
