module keyboard_ctrl (
);

// Code that takes keyboard input and converts into data used by waveform generator

endmodule
